module tt_um_example (
    input  wire [7:0] ui_in,    // Dedicated inputs
    output wire [7:0] uo_out,   // Dedicated outputs
    input  wire [7:0] uio_in,   // IOs: Input path
    output wire [7:0] uio_out,  // IOs: Output path
    output wire [7:0] uio_oe,   // IOs: Enable path (active high: 0=input, 1=output)
    input  wire       ena,      // will go high when the design is enabled
    input  wire       clk,      // clock
    input  wire       rst_n     // reset_n - low to reset
);

    // Instance of your femto system
    femto femto_instance (
        .clk(clk),
        .resetn(rst_n),
        .spi_mosi(uo_out[0]),
        .spi_miso(ui_in[0]),
        .spi_cs_n(uo_out[1]),
        .spi_clk(uo_out[2]),
        .spi_clk_ram(uo_out[3]),
        .spi_cs_n_ram(uo_out[4]),
        .spi_miso_ram(ui_in[1]),
        .spi_mosi_ram(uo_out[5]),
        .LEDS(uo_out[6]),
        .RXD(ui_in[2]),
        .TXD(uo_out[7])
    );

    // Configure bidirectional pins as inputs
    assign uio_oe = 8'b00000000;  // All bidirectional pins as inputs
    assign uio_out = 8'b00000000; // Output values for bidirectional pins

endmodule